module font_rom(clk,addr,data_reg);
input clk;
input [10:0] addr;
output reg [7:0] data_reg;

reg [7:0] data;
always @(posedge clk)
	data_reg=data;
	

always @(addr)
	case(addr)
		//S
		11'h000 : data=  8'b11111111; //
		11'h001 : data = 8'b11111111; //	
		11'h002 : data = 8'b11000000; //
		11'h003 : data = 8'b11000000; //
		11'h004 : data = 8'b11000000; //
		11'h005:  data = 8'b11000000; //
		11'h006 : data=  8'b11000000; //
		11'h007 : data = 8'b01000000; //	
		11'h008 : data = 8'b11111111; //
		11'h009 : data = 8'b11111111; //
		11'h00a : data = 8'b00000011; //
		11'h00b:  data = 8'b00000011; //
		11'h00c : data = 8'b00000011; //
		11'h00d:  data = 8'b00000011; //
		11'h00e : data = 8'b11111111; //
		11'h00f:  data = 8'b11111111; //
		//c
		11'h010 : data=  8'b00111111; //
		11'h011 : data = 8'b11111111; //	
		11'h012 : data = 8'b11110000; //
		11'h013 : data = 8'b11100000; //
		11'h014 : data = 8'b11000000 ; //
		11'h015:  data = 8'b11000000 ; //
		11'h016 : data=  8'b11000000; //
		11'h017 : data = 8'b11000000; //	
		11'h018 : data = 8'b11000000 ; //
		11'h019 : data = 8'b11000000; //
		11'h01a : data = 8'b11000000 ; //
		11'h01b:  data = 8'b11000000 ; //
		11'h01c : data = 8'b11100000 ; //
		11'h01d:  data = 8'b11110000 ; //
		11'h01e : data = 8'b11111111 ; //
		11'h01f:  data = 8'b00111111 ; //
		//O
		11'h020 : data=  8'b00000000; //
		11'h021 : data = 8'b00000000; //	
		11'h022 : data = 8'b00011000; //
		11'h023 : data = 8'b00111100; //
		11'h024 : data = 8'b01100110; //
		11'h025:  data = 8'b11000110; //
		11'h026 : data=  8'b11000011; //
		11'h027 : data = 8'b11000011; //	
		11'h028 : data = 8'b11000011; //
		11'h029 : data = 8'b11000011; //
		11'h02a : data = 8'b11000011; //
		11'h02b:  data = 8'b01100110; //
		11'h02c : data = 8'b00111100; //
		11'h02d:  data = 8'b00011000; //
		11'h02e : data = 8'b00000000; //
		11'h02f:  data = 8'b00000000; //
		//R
		11'h030 : data =  8'b11100111; //
		11'h031 : data =  8'b11101110; //	
		11'h032 : data = 8'b11101110; //
		11'h033 : data = 8'b11111100; //
		11'h034 : data = 8'b11111100; //
		11'h035:  data = 8'b11111100; //
		11'h036 : data = 8'b11111000; //
		11'h037 : data = 8'b11100000; //	
		11'h038 : data = 8'b11100000; //
		11'h039 : data = 8'b11100000; //
		11'h03a : data = 8'b11100000; //
		11'h03b:  data = 8'b11100000; //
		11'h03c : data = 8'b11100000; //
		11'h03d:  data = 8'b11100000; //
		11'h03e : data = 8'b11100000; //
		11'h03f:  data = 8'b11100000; //	
		//e
		11'h040 : data=  8'b11111111; //
		11'h041 : data = 8'b11111111; //	
		11'h042 : data = 8'b11000111; //
		11'h043 : data = 8'b11000111; //
		11'h044 : data = 8'b11000111; //
		11'h045:  data = 8'b11000111; //
		11'h046 : data = 8'b11000111; //
		11'h047 : data = 8'b11000111; //	
		11'h048 : data = 8'b11111111; //
		11'h049 : data = 8'b11111111; //
		11'h04a : data = 8'b11000000; //
		11'h04b:  data = 8'b11000000; //
		11'h04c : data = 8'b11000000; //
		11'h04d:  data = 8'b11000000; //
		11'h04e : data = 8'b11111111; //
		11'h04f:  data = 8'b11111111; //	
		//:
		11'h050 : data=  8'b00011100; //
		11'h051 : data=  8'b00011100; //	
		11'h052 : data = 8'b00011100; //
		11'h053 : data = 8'b00011100; //
		11'h054 : data = 8'b00011100; //
		11'h055:  data = 8'b00011100; //
		11'h056 : data=  8'b00000000; //
		11'h057 : data = 8'b00000000; //	
		11'h058 : data = 8'b00000000; //
		11'h059 : data = 8'b00000000; //
		11'h05a : data = 8'b00011100; //
		11'h05b:  data = 8'b00011100; //
		11'h05c : data = 8'b00011100; //
		11'h05d:  data = 8'b00011100; //
		11'h05e : data = 8'b00011100; //
		11'h05f:  data = 8'b00011100; //
		// 
		11'h060 : data=  8'b01111000; //
		11'h061 : data = 8'b11111000; //	
		11'h062 : data = 8'b11111000; //
		11'h063 : data = 8'b00111000; //
		11'h064 : data = 8'b00111000; //
		11'h065:  data = 8'b00111000; //
		11'h066 : data=  8'b00111000; //
		11'h067 : data = 8'b00111000; //	
		11'h068 : data = 8'b00111000; //
		11'h069 : data = 8'b00111000; //
		11'h06a : data = 8'b00111000; //
		11'h06b:  data = 8'b00111000; //
		11'h06c : data = 8'b00111000; //
		11'h06d:  data = 8'b00111000; //
		11'h06e : data = 8'b11111111; //
		11'h06f:  data = 8'b11111111; //
		// 
		11'h070 : data=  8'b11111111; //
		11'h071 : data = 8'b11111111 ;//	
		11'h072 : data = 8'b00000011; //
		11'h073 : data = 8'b00000011; //
		11'h074 : data = 8'b00000110; //
		11'h075:  data = 8'b00001100; //
		11'h076 : data=  8'b00011000; //
		11'h077 : data = 8'b00011000; //	
		11'h078 : data = 8'b00011000; //
		11'h079 : data = 8'b00011000; //
		11'h07a : data = 8'b00011000; //
		11'h07b:  data = 8'b00110000; //
		11'h07c : data = 8'b01100000; //
		11'h07d:  data = 8'b11000000; //
		11'h07e : data = 8'b11111111; //
		11'h07f:  data = 8'b11111111; //
		// 
		11'h080 : data=  8'b00000000; //
		11'h081 : data = 8'b00000000; //	
		11'h082 : data = 8'b00000000; //
		11'h083 : data = 8'b00000000; //
		11'h084 : data = 8'b00000000; //
		11'h085:  data = 8'b00000000; //
		11'h086 : data=  8'b00000000; //
		11'h087 : data = 8'b00000000; //	
		11'h088 : data = 8'b00000000; //
		11'h089 : data = 8'b00000000; //
		11'h08a : data = 8'b00000000; //
		11'h08b:  data = 8'b00000000; //
		11'h08c : data = 8'b00000000; //
		11'h08d:  data = 8'b00000000; //
		11'h08e : data = 8'b00000000; //
		11'h08f:  data = 8'b00000000; //
		// 
		11'h090 : data=  8'b00000000; //
		11'h091 : data = 8'b00000000; //	
		11'h092 : data = 8'b00000000; //
		11'h093 : data = 8'b00000000; //
		11'h094 : data = 8'b00000000; //
		11'h095:  data = 8'b00000000; //
		11'h096 : data=  8'b00000000; //
		11'h097 : data = 8'b00000000; //	
		11'h098 : data = 8'b00000000; //
		11'h099 : data = 8'b00000000; //
		11'h09a : data = 8'b00000000; //
		11'h09b:  data = 8'b00000000; //
		11'h09c : data = 8'b00000000; //
		11'h09d:  data = 8'b00000000; //
		11'h09e : data = 8'b00000000; //
		11'h09f:  data = 8'b00000000; //
		// B
		11'h0a0 : data=  8'b11111100; //
		11'h0a1 : data = 8'b11111110; //	
		11'h0a2 : data = 8'b11000111; //
		11'h0a3 : data = 8'b11000111; //
		11'h0a4 : data = 8'b11000111; //
		11'h0a5:  data = 8'b11000111; //
		11'h0a6 : data=  8'b11111111; //
		11'h0a7 : data = 8'b11111111; //	
		11'h0a8 : data = 8'b11111111; //
		11'h0a9 : data = 8'b11111111; //
		11'h0aa : data = 8'b11000111; //
		11'h0ab:  data = 8'b11000111; //
		11'h0ac : data = 8'b11000111; //
		11'h0ad:  data = 8'b11000111; //
		11'h0ae : data = 8'b11111110; //
		11'h0af:  data = 8'b11111100; //	
		//a
		11'h0b0 : data=  8'b00000000; //
		11'h0b1 : data = 8'b00000000; //	
		11'h0b2 : data = 8'b00000000; //
		11'h0b3 : data = 8'b11000000; //
		11'h0b4 : data = 8'b01100000; //
		11'h0b5:  data = 8'b00110000; //
		11'h0b6 : data=  8'b11110000; //
		11'h0b7 : data = 8'b11111100; //	
		11'h0b8 : data = 8'b11000110; //
		11'h0b9 : data = 8'b11000011; //
		11'h0ba : data = 8'b11000011; //
		11'h0bb:  data = 8'b11000011; //
		11'h0bc : data = 8'b11000011; //
		11'h0bd : data = 8'b11111111; //
		11'h0be : data = 8'b11111111; //
		11'h0bf:  data = 8'b00000011; //	
		// l
		11'h0c0 : data=  8'b11100000; //
		11'h0c1 : data = 8'b11100000; //	
		11'h0c2 : data = 8'b11100000; //
		11'h0c3 : data = 8'b11100000; //
		11'h0c4 : data = 8'b11100000; //
		11'h0c5:  data = 8'b11100000; //
		11'h0c6 : data=  8'b11100000; //
		11'h0c7 : data = 8'b11100000; //	
		11'h0c8 : data = 8'b11100000; //
		11'h0c9 : data = 8'b11100000; //
		11'h0ca : data = 8'b11100000; //
		11'h0cb:  data = 8'b11100000; //
		11'h0cc : data = 8'b11100000; //
		11'h0cd:  data = 8'b11100000; //
		11'h0ce : data = 8'b11111111; //
		11'h0cf:  data = 8'b11111111; //
		//l 
		11'h0d0 : data=  8'b11100000; //
		11'h0d1 : data = 8'b11100000; //	
		11'h0d2 : data = 8'b11100000; //
		11'h0d3 : data = 8'b11100000; //
		11'h0d4 : data = 8'b11100000; //
		11'h0d5:  data = 8'b11100000; //
		11'h0d6 : data=  8'b11100000; //
		11'h0d7 : data = 8'b11100000; //	
		11'h0d8 : data = 8'b11100000; //
		11'h0d9 : data = 8'b11100000; //
		11'h0da : data = 8'b11100000; //
		11'h0db:  data = 8'b11100000; //
		11'h0dc : data = 8'b11100000; //
		11'h0dd:  data = 8'b11100000; //
		11'h0de : data = 8'b11111111; //	
		//:
		11'h0e0 : data=  8'b00011100; //
		11'h0e1 : data=  8'b00011100; //	
		11'h0e2 : data = 8'b00011100; //
		11'h0e3 : data = 8'b00011100; //
		11'h0e4 : data = 8'b00011100; //
		11'h0e5:  data = 8'b00011100; //
		11'h0e6 : data = 8'b00000000; //
		11'h0e7 : data = 8'b00000000; //	
		11'h0e8 : data = 8'b00000000; //
		11'h0e9 : data = 8'b00000000; //
		11'h0ea : data = 8'b00011100; //
		11'h0eb : data = 8'b00011100; //
		11'h0ec : data = 8'b00011100; //
		11'h0ed : data = 8'b00011100; //
		11'h0ee : data = 8'b00011100; //
		11'h0ef : data = 8'b00011100; //
		// PONG 		
		//p 
		11'h100 : data=  8'b11110000; //
		11'h101 : data = 8'b11001100; //	
		11'h102 : data = 8'b11000110; //
		11'h103 : data = 8'b11000011; //
		11'h104 : data = 8'b11000011; //
		11'h105:  data = 8'b11000011; //
		11'h106 : data=  8'b11000110; //
		11'h107 : data = 8'b11001100; //	
		11'h108 : data = 8'b11011000; //
		11'h109 : data = 8'b11000000; //
		11'h10a : data = 8'b11000000; //
		11'h10b:  data = 8'b11000000; //
		11'h10c : data = 8'b11000000; //
		11'h10d:  data = 8'b11000000; //
		11'h10e : data = 8'b11000000; //
		11'h10f:  data = 8'b11000000; //
		//O
		11'h110 : data=  8'b00000000; //
		11'h111 : data = 8'b00000000; //	
		11'h112 : data = 8'b00011000; //
		11'h113 : data = 8'b00111100; //
		11'h114 : data = 8'b01100110; //
		11'h115:  data = 8'b11000110; //
		11'h116 : data=  8'b11000011; //
		11'h117 : data = 8'b11000011; //	
		11'h118 : data = 8'b11000011; //
		11'h119 : data = 8'b11000011; //
		11'h11a : data = 8'b11000011; //
		11'h11b:  data = 8'b01100110; //
		11'h11c : data = 8'b00111100; //
		11'h11d:  data = 8'b00011000; //
		11'h11e : data = 8'b00000000; //
		11'h11f:  data = 8'b00000000; //
			//n 
		11'h120 : data=  8'b00000000; //
		11'h121 : data = 8'b00000000; //	
		11'h122 : data = 8'b00000000; //
		11'h123 : data = 8'b00000000; //
		11'h124 : data = 8'b00000000; //
		11'h125:  data = 8'b00000000; //
		11'h126 : data=  8'b11111111; //
		11'h127 : data = 8'b11000111; //	
		11'h128 : data = 8'b11000011; //
		11'h129 : data = 8'b11000011; //
		11'h12a : data = 8'b11000011; //
		11'h12b:  data = 8'b11000011; //
		11'h12c : data = 8'b11000011; //
		11'h12d:  data = 8'b11000011; //
		11'h12e : data = 8'b11000011; //
		11'h12f:  data = 8'b11000011; //
		//g
		11'h130 : data=  8'b00000000; // 
		11'h131 : data = 8'b00000000; //	
		11'h132 : data = 8'b00000000; //
		11'h133 : data = 8'b00000000; //
		11'h134 : data = 8'b00000000; //
		11'h135:  data = 8'b00111111; //
		11'h136 : data=  8'b01100011; //
		11'h137 : data = 8'b11000011; //	
		11'h138 : data = 8'b11000011; //
		11'h139 : data = 8'b01100011; //
		11'h13a : data = 8'b00110011; //
		11'h13b:  data = 8'b00000011; //
		11'h13c : data = 8'b00000011; //
		11'h13d:  data = 8'b00000011; //
		11'h13e : data = 8'b11111111; //
		11'h13f:  data = 8'b11111111; //
	endcase
endmodule 